library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity memory is
Port ( address : in std_logic_vector(31 downto 0);
       write_data : in std_logic_vector(31 downto 0);
       clock : in std_logic;
       MemWrite : in std_logic;
       MemRead : in std_logic;
       read_data : out std_logic_vector(31 downto 0));
end memory;

architecture Behavioral of memory is
type mem_array is array(0 to 511) of std_logic_vector(31 downto 0);
constant gate_delay: Time := 1 ns;
begin
 mem_process: process(address, write_data, clock)
    variable data_mem : mem_array := (
    
      "00000000000000000000000000100110", -- 0
      "00000000000000000000000000100111", -- 1                                                            
      "00000000000000000000000000101000", -- 2
      "00000000000000000000000000101001", -- 3
      "00000000000000000000000000101010", -- 4       
      "00000000000000000000000000101011", -- 5 
      "00000000000000000000000000101100", -- 6
      "00000000000000000000000000101101", -- 7
      "00000000000000000000000000101110", -- 8                                                             
      "00000000000000000000000000101111", -- 9
      "00000000000000000000000000110000", -- a
      "00000000000000000000000000110001", -- b
      "00000000000000000000000000110010", -- c
      "00000000000000000000000000110011", -- d
      "00000000000000000000000000110100", -- e
      "00000000000000000000000000110101", -- f
      -- 01
      "00000000000000000000000000110110", -- 0
      "00000000000000000000000000110111", -- 1
      "00000000000000000000000000111000", -- 2
      "00000000000000000000000000111001", -- 3
      "00000000000000000000000000111010", -- 4
      "00000000000000000000000000111011",-- 5
      "00000000000000000000000000111100", -- 6
      "00000000000000000000000000111101", -- 7
      "00000000000000000000000000111110", -- 8
      "00000000000000000000000000111111", -- 9
      "00000000000000000000000001000000", -- a
      "00000000000000000000000001000001", -- b
      "00000000000000000000000001000010", -- c
      "00000000000000000000000001000011",-- d
      "00000000000000000000000001000100", -- e
      "00000000000000000000000001000101", -- f
      -- 02
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000",-- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000",-- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 03
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000",-- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 04
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000",-- a
      "00000000000000000000000000000000",-- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 05
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000",-- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000",-- f
      -- 06
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 07
      "00000000000000000000000000000000",-- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 08
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 09
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000",-- 1
      "00000000000000000000000000000000",-- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000",-- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 0a
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000",-- 9
      "00000000000000000000000000000000",-- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000",-- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 0b
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 0c
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000",-- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 0d
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 0e
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 0f
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 10
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 11
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 12
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 13
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 14
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 15
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 16
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 17
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 18
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 19
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 1a
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 1b
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 1c
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 1d
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 1e
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000", -- f
      -- 1f
      "00000000000000000000000000000000", -- 0
      "00000000000000000000000000000000", -- 1
      "00000000000000000000000000000000", -- 2
      "00000000000000000000000000000000", -- 3
      "00000000000000000000000000000000", -- 4
      "00000000000000000000000000000000", -- 5
      "00000000000000000000000000000000", -- 6
      "00000000000000000000000000000000", -- 7
      "00000000000000000000000000000000", -- 8
      "00000000000000000000000000000000", -- 9
      "00000000000000000000000000000000", -- a
      "00000000000000000000000000000000", -- b
      "00000000000000000000000000000000", -- c
      "00000000000000000000000000000000", -- d
      "00000000000000000000000000000000", -- e
      "00000000000000000000000000000000"  -- f
    );
variable addr:integer;
    begin -- the following type conversion function is in std_logic_arith
addr:=conv_integer(unsigned(address(2 downto 0)));
if MemWrite ='1' then
data_mem(addr):= write_data;
elsif MemRead='1' then
read_data <= data_mem(addr) after 10 ns;
end if;
end process;
end Behavioral;