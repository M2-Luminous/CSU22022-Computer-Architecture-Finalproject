library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity control_memory is
Port (FL : out std_logic; -- 0
    RZ : out std_logic; -- 1
    RN : out std_logic; -- 2
    RC : out std_logic; -- 3
    RV : out std_logic; -- 4
    MW : out std_logic; -- 5
    MM : out std_logic; -- 6
    RW : out std_logic; -- 7
    MD : out std_logic; -- 8
    FS : out std_logic_vector(4 downto 0); -- 9 to 13
    MB : out std_logic; -- 14
    TB : out std_logic; -- 15
    TA : out std_logic; -- 16
    TD : out std_logic; -- 17
    PL : out std_logic; -- 18
    PI : out std_logic; -- 19
    IL : out std_logic; -- 20
    MC : out std_logic; -- 21
    MS : out std_logic_vector(2 downto 0); -- 22 to 24
    NA : out std_logic_vector(16 downto 0); -- 25 to 41
    IN_CAR : in std_logic_vector(16 downto 0));
end control_memory;

architecture Behavioral of control_memory is
type mem_array is array(0 to 255) of std_logic_vector(41 downto 0);

begin
  memory_m: process(in_car)
    variable control_mem : mem_array := (
    
       "000000000000000000000000000000000000100110", -- 0 - adi dr sa const_b
       "000000000000000000000000000000000000100111", -- 1 - ld dr [sa]
       "000000000000000000000000000000000000101000", -- 2 - st [sa] sb
       "000000000000000000000000000000000000101001", -- 3 - inc dr sa
       "000000000000000000000000000000000000101010", -- 4 - not dr sa
       "000000000000000000000000000000000000101011", -- 5 - add dr sa sb
       "000000000000000000000000000000000000101100", -- 6 - b displacement
       "000000000000000000000000000000000000101101", -- 7 - bne displacement sb 
       "000000000000000000000000000000000000101110", -- 8 - nop
       "000000000000000000000000000000000000101111", -- 9 - sr dr sb
       "000000000000000000000000000000000000110000", -- a - dec dr sa
       "000000000000000000000000000000000000110001", -- b
       "000000000000000000000000000000000000110010", -- c
       "000000000000000000000000000000000000110011", -- d
       "000000000000000000000000000000000000110100", -- e
       "000000000000000000000000000000000000110101", -- f
      -- 1
       "000000000000000000000000000000000000110110", -- 0
       "000000000000000000000000000000000000110111", -- 1
       "000000000000000000000000000000000000111000", -- 2
       "000000000000000000000000000000000000111001", -- 3
       "000000000000000000000000000000000000111010", -- 4
       "000000000000000000000000000000000000111011", -- 5
       "000000000000000000000000000000000000111100", -- 6
       "000000000000000000000000000000000000111101", -- 7
       "000000000000000000000000000000000000111110", -- 8
       "000000000000000000000000000000000000111111", -- 9
       "000000000000000000000000000000000001000000", -- a
       "000000000000000000000000000000000001000001", -- b
       "000000000000000000000000000000000001000010", -- c
       "000000000000000000000000000000000001000000", -- d
       "000000000000000000000000000000000001000001", -- e
       "000000000000000000000000000000000001000010", -- f
      -- 2
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- 3
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- 4
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- 5
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- 6
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- 7
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- 8
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- 9
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- a
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- b
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- c
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- d
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- e
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000", -- f
      -- f
       "000000000000000000000000000000000000000000", -- 0
       "000000000000000000000000000000000000000000", -- 1
       "000000000000000000000000000000000000000000", -- 2
       "000000000000000000000000000000000000000000", -- 3
       "000000000000000000000000000000000000000000", -- 4
       "000000000000000000000000000000000000000000", -- 5
       "000000000000000000000000000000000000000000", -- 6
       "000000000000000000000000000000000000000000", -- 7
       "000000000000000000000000000000000000000000", -- 8
       "000000000000000000000000000000000000000000", -- 9
       "000000000000000000000000000000000000000000", -- a
       "000000000000000000000000000000000000000000", -- b
       "000000000000000000000000000000000000000000", -- c
       "000000000000000000000000000000000000000000", -- d
       "000000000000000000000000000000000000000000", -- e
       "000000000000000000000000000000000000000000"  -- f
 );
    variable addr: integer;
    variable control_out: std_logic_vector(41 downto 0);
  begin
    addr := conv_integer(IN_CAR);
    control_out := control_mem(addr);
    FL <= control_out(0);
    RZ <= control_out(1);
    RN <= control_out(2);
    RC <= control_out(3);
    RV <= control_out(4);
    MW <= control_out(5);
    MM <= control_out(6);
    RW <= control_out(7);
    MD <= control_out(8);
    FS <= control_out(13 downto 9);
    MB <= control_out(14);
    TB <= control_out(15);
    TA <= control_out(16);
    TD <= control_out(12);
    PL <= control_out(17);
    PI <= control_out(19);
    IL <= control_out(20);
    MC <= control_out(21);
    MS <= control_out(24 downto 22);
    NA <= control_out(41 downto 25);
  end process;
end Behavioral;